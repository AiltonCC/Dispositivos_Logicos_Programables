library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity TecladoSPI is
    Port ( ST : in  STD_LOGIC;
           RST : in  STD_LOGIC;
           CLK : in  STD_LOGIC;
           SS : out  STD_LOGIC;
           MISO : in  STD_LOGIC;
           SCL : out  STD_LOGIC;
           LED_SCL : out  STD_LOGIC;
           LED_SS : out  STD_LOGIC;
           SEG : out  STD_LOGIC_VECTOR (7 downto 0);
           AN : out  STD_LOGIC_VECTOR (3 downto 0));
end TecladoSPI;

architecture Behavioral of TecladoSPI is
--TECLAS
SIGNAL TECLAS: STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL SELECTOR: STD_LOGIC;

--BOTONES
--SIGNAL ST_OK: STD_LOGIC;
--SIGNAL ST_AN:  STD_LOGIC;

--OBJETO ANTI-REBOTE
--ANTIREBOTE
SIGNAL T_ESTABLE	:	INTEGER RANGE 0 TO 500_000;
SIGNAL ST_OKAN	:	STD_LOGIC;
SIGNAL ST_OK: STD_LOGIC;
SIGNAL ST_AN:  STD_LOGIC;
--DESPLIEGUE
SIGNAL DFREQ: INTEGER RANGE 0 TO 50000;
SIGNAL SEL:INTEGER RANGE 0 TO 3;
SIGNAL MUX: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL NREG: INTEGER RANGE 0 TO 15;

--COMUNICACION SPI
SIGNAL CLK_SPI, CLK_SPI_AN: STD_LOGIC;
SIGNAL CTN_CLK_SPI: INTEGER RANGE 0 TO 195;
SIGNAL INI_SPI: STD_LOGIC:='0';
SIGNAL DATO_RX: STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL NBIT: INTEGER RANGE 0  TO 16;

begin
ST_AN <= ST WHEN RISING_EDGE(CLK);
T_ESTABLE <= 0 WHEN (ST_AN = '0' AND ST = '1') OR (ST_AN = '1' AND ST = '0') OR RST = '1' OR T_ESTABLE = 500_000
					ELSE T_ESTABLE +1 WHEN RISING_EDGE(CLK);
ST_OK <= ST WHEN T_ESTABLE = 499_999 AND RISING_EDGE(CLK);
ST_OKAN <= ST_OK WHEN RISING_EDGE(CLK);
--BOTONES FLANCOS
--ST_AN <= ST_OK WHEN RISING_EDGE(CLK);

--COMUNICACION SPI
CTN_CLK_SPI <= 0 WHEN INI_SPI='0' OR CTN_CLK_SPI=195 ELSE
					CTN_CLK_SPI + 1 WHEN RISING_EDGE (CLK);
					
INI_SPI <= '0' WHEN RST='1' OR NBIT=16 ELSE 
				'1' WHEN ST_OKAN='0' AND ST_OK='1' AND RISING_EDGE(CLK);

CLK_SPI <= '0' WHEN CTN_CLK_SPI <= 97 ELSE '1';

NBIT <= 0 WHEN INI_SPI = '0' OR RST='1' ELSE
		NBIT+1 WHEN CLK_SPI_AN='1' AND CLK_SPI='0' AND RISING_EDGE(CLK);
		
SCL <= CLK_SPI;
LED_SCL <=CLK_SPI;

--FLANCO
CLK_SPI_AN <= CLK_SPI WHEN RISING_EDGE(CLK);

--SS
SS<= NOT INI_SPI;
LED_SS<= NOT INI_SPI;

PROCESS(CLK, INI_SPI, RST)

BEGIN

	IF RST='1' THEN
	DATO_RX<= X"0000";
	
	ELSIF  INI_SPI='1' AND RISING_EDGE(CLK) THEN 
	
		IF CLK_SPI_AN='1' AND CLK_SPI='0' THEN --FLANCO NEGATIVO
		DATO_RX(15 DOWNTO 1)<= DATO_RX(14 DOWNTO 0);
		DATO_RX(0) <= MISO;
		END IF;
		
	END IF;


END PROCESS;

--DESPLIEGUE
DFREQ <= 0 WHEN DFREQ=50000 ELSE
		DFREQ+1 WHEN RISING_EDGE(CLK);
		
SEL<= SEL+1 WHEN DFREQ=49999 AND RISING_EDGE(CLK);

AN<=	"0001" WHEN SEL = 0 ELSE
		"0010" WHEN SEL = 1 ELSE
		"0100" WHEN SEL = 2 ELSE
		"1000" ;
		
SEG<= X"3F" WHEN MUX = X"0" ELSE
		X"06" WHEN MUX = X"1" ELSE
		X"5B" WHEN MUX = X"2" else
		X"4F" WHEN MUX = X"3" ELSE
		X"66" WHEN MUX = X"4" ELSE
		X"6D" WHEN MUX = X"5" ELSE
		X"7D" WHEN MUX = X"6" ELSE
		X"07" WHEN MUX = X"7" ELSE
		X"7F" WHEN MUX = X"8" ELSE
		X"6F" WHEN MUX = X"9" ELSE
		X"77" WHEN MUX = X"A" ELSE
		X"7C" WHEN MUX = X"B" ELSE
		X"39" WHEN MUX = X"C" ELSE
		X"5E" WHEN MUX = X"D" ELSE
		X"79" WHEN MUX = X"E" ELSE
		X"71" ;
		
MUX <= DATO_RX (3 DOWNTO 0) WHEN SEL = 0 ELSE
		 DATO_RX (7 DOWNTO 4) WHEN SEL = 1 ELSE
		 DATO_RX (11 DOWNTO 8) WHEN SEL = 2 ELSE
		 DATO_RX (15 DOWNTO 12) ;
		 
-- CONECTAR  OBEJTO ANTI-REBOTE

end Behavioral;

