library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ComTX IS
	PORT(	DATO	:	IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			ST		:	IN STD_LOGIC;
			CLK	:	IN STD_LOGIC;
			RST	:	IN	STD_LOGIC;
			TX		:	OUT STD_LOGIC);
END ComTX;

ARCHITECTURE BEHAVIORAL OF ComTX IS
--VARIABLES PARA LA COMINICACION
SIGNAL BITRATE_TX	:	INTEGER :=0;
SIGNAL NBIT	:	INTEGER :=0;
SIGNAL INI_TX	:	STD_LOGIC;
--VARIABLES PARA ANTIREBOTE
SIGNAL T_ESTABLE	:	INTEGER RANGE 0 TO 500_000;
SIGNAL ST_AN	:	STD_LOGIC;
SIGNAL ST_OK	:	STD_LOGIC;
SIGNAL ST_ONAN	:	STD_LOGIC;
BEGIN

--ANTIREBOTE
ST_AN <= ST WHEN RISING_EDGE(CLK);
T_ESTABLE <= 0 WHEN (ST_AN = '0' AND ST = '1') OR (ST_AN = '1' AND ST = '0') OR RST = '1' OR T_ESTABLE = 500_000
					ELSE T_ESTABLE +1 WHEN RISING_EDGE(CLK);
ST_OK <= ST WHEN T_ESTABLE = 499_999 AND RISING_EDGE(CLK);
ST_ONAN <= ST_OK WHEN RISING_EDGE(CLK);

--COMUNICACION
BITRATE_TX <= 0 WHEN INI_TX = '0' OR BITRATE_TX = 5208 OR RST = '1' ELSE BITRATE_TX +1 WHEN RISING_EDGE(CLK);
NBIT <= 0 WHEN INI_TX = '0' OR RST = '1' ELSE NBIT +1 WHEN BITRATE_TX = 5207 AND RISING_EDGE(CLK);
INI_TX <= '0' WHEN RST = '1' OR NBIT = 9 ELSE '1' WHEN ST_ONAN = '0' AND ST_OK =  '1' AND RISING_EDGE(CLK);
TX <=	'1' WHEN INI_TX = '0' ELSE
		'0' WHEN NBIT = 0 ELSE
		DATO(0) WHEN NBIT = 1 ELSE
		DATO(1) WHEN NBIT = 2 ELSE
		DATO(2) WHEN NBIT = 3 ELSE
		DATO(3) WHEN NBIT = 4 ELSE
		DATO(4) WHEN NBIT = 5 ELSE
		DATO(5) WHEN NBIT = 6 ELSE
		DATO(6) WHEN NBIT = 7 ELSE
		DATO(7) WHEN NBIT = 8 ELSE
		'1';
END BEHAVIORAL;